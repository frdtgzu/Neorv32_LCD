library ieee;
use ieee.std_logic_1164.all;

library surf;
use surf.StdRtlPkg.all;
use surf.AxiStreamPkg.all;
use surf.AxiLitePkg.all;

package LcdPkg is
    
   record LcdStat

    
end package LcdPkg;

package body LcdPkg is
    
end package body LcdPkg;